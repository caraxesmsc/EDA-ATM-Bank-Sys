module ATM(
    input CLK
)